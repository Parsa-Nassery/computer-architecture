//Controller Verilog
module Controller(input clk, rst, Start, Cout1, Cout2, output reg [15:0] m, output reg Ready, en_x2, en_xx, en_xy, en_x, en_y, en_x_y, en_b0, en_b1, en_err, ld_1, ld_2, cnt1, cnt2);
	reg [3:0] nstate, pstate;
	
	parameter [3:0] idle = 0, read = 1, cal = 2, mult1 = 3, div1 = 4, sub1 = 5, div2 = 6, mult2 = 7, sub2 = 8, div3 = 9, err_init = 10, err = 11, final_err = 12, finish = 13;
	always @(pstate, Start, Cout1, Cout2) begin
		nstate = 0;
		m = 16'b0; Ready = 1'b0; en_x2 = 1'b0; en_xx = 1'b0; en_xy = 1'b0; en_x = 1'b0; en_y = 1'b0; en_x_y = 1'b0; en_b0 = 1'b0; en_b1 = 1'b0; en_err = 1'b0; ld_1 = 1'b0; ld_2 = 1'b0; cnt1 = 1'b0; cnt2 = 1'b0;
		case(pstate)
			idle: begin nstate = Start ? read : idle; Ready = 1'b1; end
			read: begin nstate = cal; ld_1 = 1'b1; ld_2 = 1'b1; end
			cal: begin nstate = Cout1 ? mult1 : cal; cnt1 = 1'b1; en_x = 1'b1; en_y = 1'b1; en_xy = 1'b1; en_xx = 1'b1; m[10] = 1'b1; m[8] = 1'd1; m[4] = 1'b1; m[2] = 1'b1; end
			mult1: begin nstate = div1; cnt2 = 1'b1; en_x2 = 1'b1; en_x_y = 1'b1; m[3] = 1'b1; m[7] = 1'b1; m[9] = 1'b1; ld_1 = 1'b1; end
			div1: begin nstate = sub1; cnt2 = 1'b1; en_x2 = 1'b1; en_x_y = 1'b1; m[15] = 1'b1; m[5] = 1'b1; end
			sub1: begin nstate = div2; cnt2 = 1'b1; en_xx = 1'b1; en_xy = 1'b1; m[13] = 1'b1; m[12] = 1'b1; end
			div2: begin nstate = mult2; cnt2 =1'b1; en_b1 = 1'b1; m[14] = 1'b1; end
			mult2: begin nstate = sub2; cnt2 = 1'b1; en_b0 = 1'b1; m[1] = 1'b1; m[3] = 1'b1; m[6] = 1'b1; m[11] = 1'b1; end
			sub2: begin nstate = div3; cnt2 = 1'b1; en_b0 = 1'b1; end
			div3: begin nstate = err_init; cnt2 = 1'b1; en_b0 = 1'b1; m[11] = 1'b1; ld_1 = 1'b1; end
			err_init: begin nstate = Cout2 ? err : err_init; cnt2 = 1'b1; end
			err: begin nstate = Cout1 ? final_err : err; cnt1 = 1'b1; en_err = 1'b1; end
			final_err: begin nstate = idle; en_err = 1'b1; end
			default: nstate = idle;
		endcase
	end
	always @(posedge clk, posedge rst) begin
		if(rst)
			pstate <= idle;
		else
			pstate <= nstate;
	end
endmodule		 
